module TestMyBundle(
  input   clock,
  input   reset
);
endmodule
